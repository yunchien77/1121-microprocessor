




		
		
		
		
		
		
		
		
		
		
		
		