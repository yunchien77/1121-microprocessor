LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY SevenSegment is
	PORT ( Z0, Y0, X0, W0, Z1, Y1, X1, W1: IN std_logic;
			 a0, b0, c0, d0, e0, f0, g0, a1, b1, c1, d1, e1, f1, g1: OUT std_logic);
END SevenSegment;

ARCHITECTURE func of SevenSegment is
BEGIN
	a0 <= (NOT W0 AND NOT X0 AND NOT Y0 AND Z0) 
			OR (NOT W0 AND X0 AND NOT Y0 AND NOT Z0) 
			OR (W0 AND NOT X0 AND Y0 AND Z0) 
			OR (W0 AND X0 AND NOT Y0);
	b0 <= (NOT W0 AND X0 AND NOT Y0 AND Z0) 
			OR (NOT W0 AND X0 AND Y0 AND NOT Z0)
			OR (W0 AND NOT X0 AND Y0 AND Z0)
			OR (W0 AND X0 AND NOT Z0)
			OR (W0 AND X0 AND Y0);
	c0 <= (NOT W0 AND NOT X0 AND Y0 AND NOT Z0)
			OR (W0 AND X0 AND NOT Z0)
			OR (W0 AND X0 AND Y0);
	d0 <= (NOT X0 AND NOT Y0 AND Z0)
			OR (NOT W0 AND X0 AND NOT Y0 AND NOT Z0)
			OR (X0 AND Y0 AND Z0)
			OR (W0 AND NOT X0 AND Y0 AND NOT Z0);
	e0 <= (NOT W0 AND Z0) 
			OR (NOT W0 AND X0 AND NOT Y0)
			OR (NOT X0 AND NOT Y0 AND Z0);
	f0 <= (NOT W0 AND NOT X0 AND Z0)
			OR (NOT W0 AND NOT X0 AND Y0)
			OR (NOT W0 AND Y0 AND Z0)
			OR (W0 AND X0 AND NOT Y0);
	g0 <= (NOT W0 AND NOT X0 AND NOT Y0)
			OR (NOT W0 AND X0 AND Y0 AND Z0);
			
	a1 <= (NOT W1 AND NOT X1 AND NOT Y1 AND Z1) 
			OR (NOT W1 AND X1 AND NOT Y1 AND NOT Z1) 
			OR (W1 AND NOT X1 AND Y1 AND Z1) 
			OR (W1 AND X1 AND NOT Y1);
	b1 <= (NOT W1 AND X1 AND NOT Y1 AND Z1) 
			OR (NOT W1 AND X1 AND Y1 AND NOT Z1)
			OR (W1 AND NOT X1 AND Y1 AND Z1)
			OR (W1 AND X1 AND NOT Z1)
			OR (W1 AND X1 AND Y1);
	c1 <= (NOT W1 AND NOT X1 AND Y1 AND NOT Z1)
			OR (W1 AND X1 AND NOT Z1)
			OR (W1 AND X1 AND Y1);
	d1 <= (NOT X1 AND NOT Y1 AND Z1)
			OR (NOT W1 AND X1 AND NOT Y1 AND NOT Z1)
			OR (X1 AND Y1 AND Z1)
			OR (W1 AND NOT X1 AND Y1 AND NOT Z1);
	e1 <= (NOT W1 AND Z1) 
			OR (NOT W1 AND X1 AND NOT Y1)
			OR (NOT X1 AND NOT Y1 AND Z1);
	f1 <= (NOT W1 AND NOT X1 AND Z1)
			OR (NOT W1 AND NOT X1 AND Y1)
			OR (NOT W1 AND Y1 AND Z1)
			OR (W1 AND X1 AND NOT Y1);
	g1 <= (NOT W1 AND NOT X1 AND NOT Y1)
			OR (NOT W1 AND X1 AND Y1 AND Z1);
END func;